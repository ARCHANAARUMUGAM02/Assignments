`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02.09.2025 10:25:54
// Design Name: 
// Module Name: fsm_one_testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fsm_one_testbench();
reg clk,rst,x;
wire y;
fsm_sequence_detector uut (.clk(clk),.rst(rst),.x(x),.y(y));
reg[15:0]test_vector;
integer i;
always#5 clk=~clk;
initial begin
        clk = 0; rst = 1; x = 0;
        #12 rst = 0;
        test_vector= 16'b0101101111010100;
        for (i = 15; i >= 0; i = i - 1) begin
            x = test_vector[i];
            #10;
        end
        #20 $finish;
    end

endmodule

