`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 25.07.2025 18:19:21
// Design Name: 
// Module Name: part_selectt
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module part_selectt();
reg[7:0]bus;
reg[3:0]out;
initial begin
bus=8'b00001111;
out=4'b1111;
end
endmodule
