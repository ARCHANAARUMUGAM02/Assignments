`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01.08.2025 18:27:03
// Design Name: 
// Module Name: rtl_snippet
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module rtl_snippet(input wire clk,input wire x1,x2,x3,output reg e,f);
wire x1,x2,x3;
assign d1=x3|f;
assign d2=x1&x2;
always@(posedge clk)begin
e<=d1;
f<=d2;
end
endmodule
