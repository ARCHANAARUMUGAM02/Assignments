`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 25.07.2025 17:37:53
// Design Name: 
// Module Name: reall_ttime
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module reall_ttime();
real delta_1,delta_2;
  integer int_value_1,int value_2;
initial begin
delta_1=4e10;
  int_value_1=delta_1;
  delta_2=2.18;
  int_value_2=delta_2;
end
endmodule
